module wlr

pub struct C.wlr_session {
}

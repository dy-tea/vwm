module xkb

pub enum Keysym as u32 {
	nosymbol    = 0x000000
	voidsymbol  = 0xffffff
	backspace   = 0xff08
	tab         = 0xff09
	linefeed    = 0xff0a
	clear       = 0xff0b
	return      = 0xff0d
	pause       = 0xff13
	scroll_lock = 0xff14
	sys_req     = 0xff15
	escape      = 0xff1b
	delete      = 0xffff

	multi_key         = 0xff20
	codeinput         = 0xff37
	singlecandidate   = 0xff3c
	multiplecandidate = 0xff3d
	previouscandidate = 0xff3e

	kanji             = 0xff21
	muhenkan          = 0xff22
	henkan            = 0xff23
	romaji            = 0xff24
	hiragana          = 0xff25
	katakana          = 0xff26
	hiragana_katakana = 0xff27
	zenkaku           = 0xff28
	hankaku           = 0xff29
	zenkaku_hankaku   = 0xff2a
	touroku           = 0xff2b
	massyo            = 0xff2c
	kana_lock         = 0xff2d
	kana_shift        = 0xff2e
	eisu_shift        = 0xff2f
	eisu_toggle       = 0xff30

	home  = 0xff50
	left  = 0xff51
	up    = 0xff52
	right = 0xff53
	down  = 0xff54
	prior = 0xff55
	next  = 0xff56
	end   = 0xff57
	begin = 0xff58

	select      = 0xff60
	print       = 0xff61
	execute     = 0xff62
	insert      = 0xff63
	undo        = 0xff65
	redo        = 0xff66
	menu        = 0xff67
	find        = 0xff68
	cancel      = 0xff69
	help        = 0xff6a
	break       = 0xff6b
	mode_switch = 0xff7e
	num_lock    = 0xff7f

	kp_space     = 0xff80
	kp_tab       = 0xff89
	kp_enter     = 0xff8d
	kp_f1        = 0xff91
	kp_f2        = 0xff92
	kp_f3        = 0xff93
	kp_f4        = 0xff94
	kp_home      = 0xff95
	kp_left      = 0xff96
	kp_up        = 0xff97
	kp_right     = 0xff98
	kp_down      = 0xff99
	kp_prior     = 0xff9a
	kp_next      = 0xff9b
	kp_end       = 0xff9c
	kp_begin     = 0xff9d
	kp_insert    = 0xff9e
	kp_delete    = 0xff9f
	kp_equal     = 0xffbd
	kp_multiply  = 0xffaa
	kp_add       = 0xffab
	kp_separator = 0xffac
	kp_subtract  = 0xffad
	kp_decimal   = 0xffae
	kp_divide    = 0xffaf

	kp_0 = 0xffb0
	kp_1 = 0xffb1
	kp_2 = 0xffb2
	kp_3 = 0xffb3
	kp_4 = 0xffb4
	kp_5 = 0xffb5
	kp_6 = 0xffb6
	kp_7 = 0xffb7
	kp_8 = 0xffb8
	kp_9 = 0xffb9

	f1  = 0xffbe
	f2  = 0xffbf
	f3  = 0xffc0
	f4  = 0xffc1
	f5  = 0xffc2
	f6  = 0xffc3
	f7  = 0xffc4
	f8  = 0xffc5
	f9  = 0xffc6
	f10 = 0xffc7
	f11 = 0xffc8
	f12 = 0xffc9
	f13 = 0xffca
	f14 = 0xffcb
	f15 = 0xffcc
	f16 = 0xffcd
	f17 = 0xffce
	f18 = 0xffcf
	f19 = 0xffd0
	f20 = 0xffd1
	f21 = 0xffd2
	f22 = 0xffd3
	f23 = 0xffd4
	f24 = 0xffd5
	f25 = 0xffd6
	f26 = 0xffd7
	f27 = 0xffd8
	f28 = 0xffd9
	f29 = 0xffda
	f30 = 0xffdb
	f31 = 0xffdc
	f32 = 0xffdd
	f33 = 0xffde
	f34 = 0xffdf
	f35 = 0xffe0

	shift_l    = 0xffe1
	shift_r    = 0xffe2
	control_l  = 0xffe3
	control_r  = 0xffe4
	caps_lock  = 0xffe5
	shift_lock = 0xffe6

	meta_l  = 0xffe7
	meta_r  = 0xffe8
	alt_l   = 0xffe9
	alt_r   = 0xffea
	super_l = 0xffeb
	super_r = 0xffec
	hyper_l = 0xffed
	hyper_r = 0xffee

	iso_lock             = 0xfe01
	iso_level2_latch     = 0xfe02
	iso_level3_shift     = 0xfe03
	iso_level3_latch     = 0xfe04
	iso_level3_lock      = 0xfe05
	iso_level5_shift     = 0xfe11
	iso_level5_latch     = 0xfe12
	iso_level5_lock      = 0xfe13
	iso_group_latch      = 0xfe06
	iso_group_lock       = 0xfe07
	iso_next_group       = 0xfe08
	iso_next_group_lock  = 0xfe09
	iso_prev_group       = 0xfe0a
	iso_prev_group_lock  = 0xfe0b
	iso_first_group      = 0xfe0c
	iso_first_group_lock = 0xfe0d
	iso_last_group       = 0xfe0e
	iso_last_group_lock  = 0xfe0f

	iso_left_tab                = 0xfe20
	iso_move_line_up            = 0xfe21
	iso_move_line_down          = 0xfe22
	iso_partial_line_up         = 0xfe23
	iso_partial_line_down       = 0xfe24
	iso_partial_space_left      = 0xfe25
	iso_partial_space_right     = 0xfe26
	iso_set_margin_left         = 0xfe27
	iso_set_margin_right        = 0xfe28
	iso_release_margin_left     = 0xfe29
	iso_release_margin_right    = 0xfe2a
	iso_release_both_margins    = 0xfe2b
	iso_fast_cursor_left        = 0xfe2c
	iso_fast_cursor_right       = 0xfe2d
	iso_fast_cursor_up          = 0xfe2e
	iso_fast_cursor_down        = 0xfe2f
	iso_continuous_underline    = 0xfe30
	iso_discontinuous_underline = 0xfe31
	iso_emphasize               = 0xfe32
	iso_center_object           = 0xfe33
	iso_enter                   = 0xfe34

	dead_grave              = 0xfe50
	dead_acute              = 0xfe51
	dead_circumflex         = 0xfe52
	dead_tilde              = 0xfe53
	dead_macron             = 0xfe54
	dead_breve              = 0xfe55
	dead_abovedot           = 0xfe56
	dead_diaeresis          = 0xfe57
	dead_abovering          = 0xfe58
	dead_doubleacute        = 0xfe59
	dead_caron              = 0xfe5a
	dead_cedilla            = 0xfe5b
	dead_ogonek             = 0xfe5c
	dead_iota               = 0xfe5d
	dead_voiced_sound       = 0xfe5e
	dead_semivoiced_sound   = 0xfe5f
	dead_belowdot           = 0xfe60
	dead_hook               = 0xfe61
	dead_horn               = 0xfe62
	dead_stroke             = 0xfe63
	dead_abovecomma         = 0xfe64
	dead_abovereversedcomma = 0xfe65
	dead_doublegrave        = 0xfe66
	dead_belowring          = 0xfe67
	dead_belowmacron        = 0xfe68
	dead_belowcircumflex    = 0xfe69
	dead_belowtilde         = 0xfe6a
	dead_belowbreve         = 0xfe6b
	dead_belowdiaeresis     = 0xfe6c
	dead_invertedbreve      = 0xfe6d
	dead_belowcomma         = 0xfe6e
	dead_currency           = 0xfe6f

	dead_lowline            = 0xfe90
	dead_aboveverticalline  = 0xfe91
	dead_belowverticalline  = 0xfe92
	dead_longsolidusoverlay = 0xfe93

	dead_a           = 0xfe80
	dead_a_upper     = 0xfe81
	dead_e           = 0xfe82
	dead_e_upper     = 0xfe83
	dead_i           = 0xfe84
	dead_i_upper     = 0xfe85
	dead_o           = 0xfe86
	dead_o_upper     = 0xfe87
	dead_u           = 0xfe88
	dead_u_upper     = 0xfe89
	dead_schwa       = 0xfe8a
	dead_schwa_upper = 0xfe8b

	dead_greek = 0xfe8c
	dead_hamza = 0xfe8d

	first_virtual_screen = 0xfed0
	prev_virtual_screen  = 0xfed1
	next_virtual_screen  = 0xfed2
	last_virtual_screen  = 0xfed4
	terminate_server     = 0xfed5

	accessx_enable          = 0xfe70
	accessx_feedback_enable = 0xfe71
	repeatkeys_enable       = 0xfe72
	slowkeys_enable         = 0xfe73
	bouncekeys_enable       = 0xfe74
	stickykeys_enable       = 0xfe75
	mousekeys_enable        = 0xfe76
	mousekeys_accel_enable  = 0xfe77
	overlay1_enable         = 0xfe78
	overlay2_enable         = 0xfe79
	audiblebell_enable      = 0xfe7a

	pointer_left          = 0xfee0
	pointer_right         = 0xfee1
	pointer_up            = 0xfee2
	pointer_down          = 0xfee3
	pointer_upleft        = 0xfee4
	pointer_upright       = 0xfee5
	pointer_downleft      = 0xfee6
	pointer_downright     = 0xfee7
	pointer_button_dflt   = 0xfee8
	pointer_button1       = 0xfee9
	pointer_button2       = 0xfeea
	pointer_button3       = 0xfeeb
	pointer_button4       = 0xfeec
	pointer_button5       = 0xfeed
	pointer_dblclick_dflt = 0xfeee
	pointer_dblclick1     = 0xfeef
	pointer_dblclick2     = 0xfef0
	pointer_dblclick3     = 0xfef1
	pointer_dblclick4     = 0xfef2
	pointer_dblclick5     = 0xfef3
	pointer_drag_dflt     = 0xfef4
	pointer_drag1         = 0xfef5
	pointer_drag2         = 0xfef6
	pointer_drag3         = 0xfef7
	pointer_drag4         = 0xfef8
	pointer_drag5         = 0xfefd

	pointer_enablekeys  = 0xfef9
	pointer_accelerate  = 0xfefa
	pointer_dfltbtnnext = 0xfefb
	pointer_dfltbtnprev = 0xfefc

	ch              = 0xfea0
	ch_upper        = 0xfea1
	ch_upper_upper  = 0xfea2
	c_h             = 0xfea3
	c_h_upper       = 0xfea4
	c_h_upper_upper = 0xfea5

	_3270_duplicate    = 0xfd01
	_3270_fieldmark    = 0xfd02
	_3270_right2       = 0xfd03
	_3270_left2        = 0xfd04
	_3270_backtab      = 0xfd05
	_3270_eraseeof     = 0xfd06
	_3270_eraseinput   = 0xfd07
	_3270_reset        = 0xfd08
	_3270_quit         = 0xfd09
	_3270_pa1          = 0xfd0a
	_3270_pa2          = 0xfd0b
	_3270_pa3          = 0xfd0c
	_3270_test         = 0xfd0d
	_3270_attn         = 0xfd0e
	_3270_cursorblink  = 0xfd0f
	_3270_altcursor    = 0xfd10
	_3270_keyclick     = 0xfd11
	_3270_jump         = 0xfd12
	_3270_ident        = 0xfd13
	_3270_rule         = 0xfd14
	_3270_copy         = 0xfd15
	_3270_play         = 0xfd16
	_3270_setup        = 0xfd17
	_3270_record       = 0xfd18
	_3270_changescreen = 0xfd19
	_3270_deleteword   = 0xfd1a
	_3270_exselect     = 0xfd1b
	_3270_cursorselect = 0xfd1c
	_3270_printscreen  = 0xfd1d
	_3270_enter        = 0xfd1e

	space        = 0x0020
	exclam       = 0x0021
	quotedbl     = 0x0022
	numbersign   = 0x0023
	dollar       = 0x0024
	percent      = 0x0025
	ampersand    = 0x0026
	apostrophe   = 0x0027
	parenleft    = 0x0028
	parenright   = 0x0029
	asterisk     = 0x002a
	plus         = 0x002b
	comma        = 0x002c
	minus        = 0x002d
	period       = 0x002e
	slash        = 0x002f
	_0           = 0x0030
	_1           = 0x0031
	_2           = 0x0032
	_3           = 0x0033
	_4           = 0x0034
	_5           = 0x0035
	_6           = 0x0036
	_7           = 0x0037
	_8           = 0x0038
	_9           = 0x0039
	colon        = 0x003a
	semicolon    = 0x003b
	less         = 0x003c
	equal        = 0x003d
	greater      = 0x003e
	question     = 0x003f
	at           = 0x0040
	a_upper      = 0x0041
	b_upper      = 0x0042
	c_upper      = 0x0043
	d_upper      = 0x0044
	e_upper      = 0x0045
	f_upper      = 0x0046
	g_upper      = 0x0047
	h_upper      = 0x0048
	i_upper      = 0x0049
	j_upper      = 0x004a
	k_upper      = 0x004b
	l_upper      = 0x004c
	m_upper      = 0x004d
	n_upper      = 0x004e
	o_upper      = 0x004f
	p_upper      = 0x0050
	q_upper      = 0x0051
	r_upper      = 0x0052
	s_upper      = 0x0053
	t_upper      = 0x0054
	u_upper      = 0x0055
	v_upper      = 0x0056
	w_upper      = 0x0057
	x_upper      = 0x0058
	y_upper      = 0x0059
	z_upper      = 0x005a
	bracketleft  = 0x005b
	backslash    = 0x005c
	bracketright = 0x005d
	asciicircum  = 0x005e
	underscore   = 0x005f
	grave        = 0x0060
	a            = 0x0061
	b            = 0x0062
	c            = 0x0063
	d            = 0x0064
	e            = 0x0065
	f            = 0x0066
	g            = 0x0067
	h            = 0x0068
	i            = 0x0069
	j            = 0x006a
	k            = 0x006b
	l            = 0x006c
	m            = 0x006d
	n            = 0x006e
	o            = 0x006f
	p            = 0x0070
	q            = 0x0071
	r            = 0x0072
	s            = 0x0073
	t            = 0x0074
	u            = 0x0075
	v            = 0x0076
	w            = 0x0077
	x            = 0x0078
	y            = 0x0079
	z            = 0x007a
	braceleft    = 0x007b
	bar          = 0x007c
	braceright   = 0x007d
	asciitilde   = 0x007e

	nobreakspace      = 0x00a0
	exclamdown        = 0x00a1
	cent              = 0x00a2
	sterling          = 0x00a3
	currency          = 0x00a4
	yen               = 0x00a5
	brokenbar         = 0x00a6
	section           = 0x00a7
	diaeresis         = 0x00a8
	copyright         = 0x00a9
	ordfeminine       = 0x00aa
	guillemetleft     = 0x00ab
	notsign           = 0x00ac
	hyphen            = 0x00ad
	registered        = 0x00ae
	macron            = 0x00af
	degree            = 0x00b0
	plusminus         = 0x00b1
	twosuperior       = 0x00b2
	threesuperior     = 0x00b3
	acute             = 0x00b4
	mu                = 0x00b5
	paragraph         = 0x00b6
	periodcentered    = 0x00b7
	cedilla           = 0x00b8
	onesuperior       = 0x00b9
	ordmasculine      = 0x00ba
	guillemetright    = 0x00bb
	onequarter        = 0x00bc
	onehalf           = 0x00bd
	threequarters     = 0x00be
	questiondown      = 0x00bf
	agrave_upper      = 0x00c0
	aacute_upper      = 0x00c1
	acircumflex_upper = 0x00c2
	atilde_upper      = 0x00c3
	adiaeresis_upper  = 0x00c4
	aring_upper       = 0x00c5
	ae_upper          = 0x00c6
	ccedilla_upper    = 0x00c7
	egrave_upper      = 0x00c8
	eacute_upper      = 0x00c9
	ecircumflex_upper = 0x00ca
	ediaeresis_upper  = 0x00cb
	igrave_upper      = 0x00cc
	iacute_upper      = 0x00cd
	icircumflex_upper = 0x00ce
	idiaeresis_upper  = 0x00cf
	eth_upper         = 0x00d0
	ntilde_upper      = 0x00d1
	ograve_upper      = 0x00d2
	oacute_upper      = 0x00d3
	ocircumflex_upper = 0x00d4
	otilde_upper      = 0x00d5
	odiaeresis_upper  = 0x00d6
	multiply          = 0x00d7
	oslash_upper      = 0x00d8
	ugrave_upper      = 0x00d9
	uacute_upper      = 0x00da
	ucircumflex_upper = 0x00db
	udiaeresis_upper  = 0x00dc
	yacute_upper      = 0x00dd
	thorn_upper       = 0x00de
	ssharp_upper      = 0x00df
	agrave            = 0x00e0
	aacute            = 0x00e1
	acircumflex       = 0x00e2
	atilde            = 0x00e3
	adiaeresis        = 0x00e4
	aring             = 0x00e5
	ae                = 0x00e6
	ccedilla          = 0x00e7
	egrave            = 0x00e8
	eacute            = 0x00e9
	ecircumflex       = 0x00ea
	ediaeresis        = 0x00eb
	igrave            = 0x00ec
	iacute            = 0x00ed
	icircumflex       = 0x00ee
	idiaeresis        = 0x00ef
	eth               = 0x00f0
	ntilde            = 0x00f1
	ograve            = 0x00f2
	oacute            = 0x00f3
	ocircumflex       = 0x00f4
	otilde            = 0x00f5
	odiaeresis        = 0x00f6
	division          = 0x00f7
	oslash            = 0x00f8
	ugrave            = 0x00f9
	uacute            = 0x00fa
	ucircumflex       = 0x00fb
	udiaeresis        = 0x00fc
	yacute            = 0x00fd
	thorn             = 0x00fe
	ydiaeresis        = 0x00ff

	aogonek_upper      = 0x01a1
	breve              = 0x01a2
	lstroke_upper      = 0x01a3
	lcaron_upper       = 0x01a5
	sacute_upper       = 0x01a6
	scaron_upper       = 0x01a9
	scedilla_upper     = 0x01aa
	tcaron_upper       = 0x01ab
	zacute_upper       = 0x01ac
	zcaron_upper       = 0x01ae
	zabovedot_upper    = 0x01af
	aogonek            = 0x01b1
	ogonek             = 0x01b2
	lstroke            = 0x01b3
	lcaron             = 0x01b5
	sacute             = 0x01b6
	caron              = 0x01b7
	scaron             = 0x01b9
	scedilla           = 0x01ba
	tcaron             = 0x01bb
	zacute             = 0x01bc
	doubleacute        = 0x01bd
	zcaron             = 0x01be
	zabovedot          = 0x01bf
	racute_upper       = 0x01c0
	abreve_upper       = 0x01c3
	lacute_upper       = 0x01c5
	cacute_upper       = 0x01c6
	ccaron_upper       = 0x01c8
	eogonek_upper      = 0x01ca
	ecaron_upper       = 0x01cc
	dcaron_upper       = 0x01cf
	dstroke_upper      = 0x01d0
	nacute_upper       = 0x01d1
	ncaron_upper       = 0x01d2
	odoubleacute_upper = 0x01d5
	rcaron_upper       = 0x01d8
	uring_upper        = 0x01d9
	udoubleacute_upper = 0x01db
	tcedilla_upper     = 0x01de
	racute             = 0x01e0
	abreve             = 0x01e3
	lacute             = 0x01e5
	cacute             = 0x01e6
	ccaron             = 0x01e8
	eogonek            = 0x01ea
	ecaron             = 0x01ec
	dcaron             = 0x01ef
	dstroke            = 0x01f0
	nacute             = 0x01f1
	ncaron             = 0x01f2
	odoubleacute       = 0x01f5
	rcaron             = 0x01f8
	uring              = 0x01f9
	udoubleacute       = 0x01fb
	tcedilla           = 0x01fe
	abovedot           = 0x01ff
	hstroke_upper      = 0x02a1
	hcircumflex_upper  = 0x02a6
	iabovedot_upper    = 0x02a9
	gbreve_upper       = 0x02ab
	jcircumflex_upper  = 0x02ac
	hstroke            = 0x02b1
	hcircumflex        = 0x02b6
	idotless           = 0x02b9
	gbreve             = 0x02bb
	jcircumflex        = 0x02bc
	cabovedot_upper    = 0x02c5
	ccircumflex_upper  = 0x02c6
	gabovedot_upper    = 0x02d5
	gcircumflex_upper  = 0x02d8
	ubreve_upper       = 0x02dd
	scircumflex_upper  = 0x02de
	cabovedot          = 0x02e5
	ccircumflex        = 0x02e6
	gabovedot          = 0x02f5
	gcircumflex        = 0x02f8
	ubreve             = 0x02fd
	scircumflex        = 0x02fe

	kra             = 0x03a2
	rcedilla_upper  = 0x03a3
	itilde_upper    = 0x03a5
	lcedilla_upper  = 0x03a6
	emacron_upper   = 0x03aa
	gcedilla_upper  = 0x03ab
	tslash_upper    = 0x03ac
	rcedilla        = 0x03b3
	itilde          = 0x03b5
	lcedilla        = 0x03b6
	emacron         = 0x03ba
	gcedilla        = 0x03bb
	tslash          = 0x03bc
	eng_upper       = 0x03bd
	eng             = 0x03bf
	amacron_upper   = 0x03c0
	iogonek_upper   = 0x03c7
	eabovedot_upper = 0x03cc
	imacron_upper   = 0x03cf
	ncedilla_upper  = 0x03d1
	omacron_upper   = 0x03d2
	kcedilla_upper  = 0x03d3
	uogonek_upper   = 0x03d9
	utilde_upper    = 0x03dd
	umacron_upper   = 0x03de
	amacron         = 0x03e0
	iogonek         = 0x03e7
	eabovedot       = 0x03ec
	imacron         = 0x03ef
	ncedilla        = 0x03f1
	omacron         = 0x03f2
	kcedilla        = 0x03f3
	uogonek         = 0x03f9
	utilde          = 0x03fd
	umacron         = 0x03fe

	wcircumflex_upper       = 0x1000174
	wcircumflex             = 0x1000175
	ycircumflex_upper       = 0x1000176
	ycircumflex             = 0x1000177
	babovedot_upper         = 0x1001e02
	babovedot               = 0x1001e03
	dabovedot_upper         = 0x1001e0a
	dabovedot               = 0x1001e0b
	fabovedot_upper         = 0x1001e1e
	fabovedot               = 0x1001e1f
	mabovedot_upper         = 0x1001e40
	mabovedot               = 0x1001e41
	pabovedot_upper         = 0x1001e56
	pabovedot               = 0x1001e57
	sabovedot_upper         = 0x1001e60
	sabovedot               = 0x1001e61
	tabovedot_upper         = 0x1001e6a
	tabovedot               = 0x1001e6b
	wgrave_upper            = 0x1001e80
	wgrave                  = 0x1001e81
	wacute_upper            = 0x1001e82
	wacute                  = 0x1001e83
	wdiaeresis_upper        = 0x1001e84
	wdiaeresis              = 0x1001e85
	ygrave_upper            = 0x1001ef2
	ygrave                  = 0x1001ef3
	oe                      = 0x13bc
	oe_upper                = 0x13bd
	ydiaeresis_upper        = 0x13be
	overline                = 0x047e
	kana_fullstop           = 0x04a1
	kana_openingbracket     = 0x04a2
	kana_closingbracket     = 0x04a3
	kana_comma              = 0x04a4
	kana_conjunctive        = 0x04a5
	kana_wo_small           = 0x04a6
	kana_a_small            = 0x04a7
	kana_i_small            = 0x04a8
	kana_u_small            = 0x04a9
	kana_e_small            = 0x04aa
	kana_o_small            = 0x04ab
	kana_ya_small           = 0x04ac
	kana_yu_small           = 0x04ad
	kana_yo_small           = 0x04ae
	kana_tsu_small          = 0x04af
	prolongedsound          = 0x04b0
	kana_a                  = 0x04b1
	kana_i                  = 0x04b2
	kana_u                  = 0x04b3
	kana_e                  = 0x04b4
	kana_o                  = 0x04b5
	kana_ka                 = 0x04b6
	kana_ki                 = 0x04b7
	kana_ku                 = 0x04b8
	kana_ke                 = 0x04b9
	kana_ko                 = 0x04ba
	kana_sa                 = 0x04bb
	kana_shi                = 0x04bc
	kana_su                 = 0x04bd
	kana_se                 = 0x04be
	kana_so                 = 0x04bf
	kana_ta                 = 0x04c0
	kana_chi                = 0x04c1
	kana_tsu                = 0x04c2
	kana_te                 = 0x04c3
	kana_to                 = 0x04c4
	kana_na                 = 0x04c5
	kana_ni                 = 0x04c6
	kana_nu                 = 0x04c7
	kana_ne                 = 0x04c8
	kana_no                 = 0x04c9
	kana_ha                 = 0x04ca
	kana_hi                 = 0x04cb
	kana_fu                 = 0x04cc
	kana_he                 = 0x04cd
	kana_ho                 = 0x04ce
	kana_ma                 = 0x04cf
	kana_mi                 = 0x04d0
	kana_mu                 = 0x04d1
	kana_me                 = 0x04d2
	kana_mo                 = 0x04d3
	kana_ya                 = 0x04d4
	kana_yu                 = 0x04d5
	kana_yo                 = 0x04d6
	kana_ra                 = 0x04d7
	kana_ri                 = 0x04d8
	kana_ru                 = 0x04d9
	kana_re                 = 0x04da
	kana_ro                 = 0x04db
	kana_wa                 = 0x04dc
	kana_n                  = 0x04dd
	voicedsound             = 0x04de
	semivoicedsound         = 0x04df
	farsi_0                 = 0x10006f0
	farsi_1                 = 0x10006f1
	farsi_2                 = 0x10006f2
	farsi_3                 = 0x10006f3
	farsi_4                 = 0x10006f4
	farsi_5                 = 0x10006f5
	farsi_6                 = 0x10006f6
	farsi_7                 = 0x10006f7
	farsi_8                 = 0x10006f8
	farsi_9                 = 0x10006f9
	arabic_percent          = 0x100066a
	arabic_superscript_alef = 0x1000670
	arabic_tteh             = 0x1000679
	arabic_peh              = 0x100067e
	arabic_tcheh            = 0x1000686
	arabic_ddal             = 0x1000688
	arabic_rreh             = 0x1000691
	arabic_comma            = 0x05ac
	arabic_fullstop         = 0x10006d4
	arabic_0                = 0x1000660
	arabic_1                = 0x1000661
	arabic_2                = 0x1000662
	arabic_3                = 0x1000663
	arabic_4                = 0x1000664
	arabic_5                = 0x1000665
	arabic_6                = 0x1000666
	arabic_7                = 0x1000667
	arabic_8                = 0x1000668
	arabic_9                = 0x1000669
	arabic_semicolon        = 0x05bb
	arabic_question_mark    = 0x05bf
	arabic_hamza            = 0x05c1
	arabic_maddaonalef      = 0x05c2
	arabic_hamzaonalef      = 0x05c3
	arabic_hamzaonwaw       = 0x05c4
	arabic_hamzaunderalef   = 0x05c5
	arabic_hamzaonyeh       = 0x05c6
	arabic_alef             = 0x05c7
	arabic_beh              = 0x05c8
	arabic_tehmarbuta       = 0x05c9
	arabic_teh              = 0x05ca
	arabic_theh             = 0x05cb
	arabic_jeem             = 0x05cc
	arabic_hah              = 0x05cd
	arabic_khah             = 0x05ce
	arabic_dal              = 0x05cf
	arabic_thal             = 0x05d0
	arabic_ra               = 0x05d1
	arabic_zain             = 0x05d2
	arabic_seen             = 0x05d3
	arabic_sheen            = 0x05d4
	arabic_sad              = 0x05d5
	arabic_dad              = 0x05d6
	arabic_tah              = 0x05d7
	arabic_zah              = 0x05d8
	arabic_ain              = 0x05d9
	arabic_ghain            = 0x05da
	arabic_tatweel          = 0x05e0
	arabic_feh              = 0x05e1
	arabic_qaf              = 0x05e2
	arabic_kaf              = 0x05e3
	arabic_lam              = 0x05e4
	arabic_meem             = 0x05e5
	arabic_noon             = 0x05e6
	arabic_ha               = 0x05e7
	arabic_waw              = 0x05e8
	arabic_alefmaksura      = 0x05e9
	arabic_yeh              = 0x05ea
	arabic_fathatan         = 0x05eb
	arabic_dammatan         = 0x05ec
	arabic_kasratan         = 0x05ed
	arabic_fatha            = 0x05ee
	arabic_damma            = 0x05ef
	arabic_kasra            = 0x05f0
	arabic_shadda           = 0x05f1
	arabic_sukun            = 0x05f2
	arabic_madda_above      = 0x1000653
	arabic_hamza_above      = 0x1000654
	arabic_hamza_below      = 0x1000655
	arabic_jeh              = 0x1000698
	arabic_veh              = 0x10006a4
	arabic_keheh            = 0x10006a9
	arabic_gaf              = 0x10006af
	arabic_noon_ghunna      = 0x10006ba
	arabic_heh_doachashmee  = 0x10006be
	farsi_yeh               = 0x10006cc
	arabic_yeh_baree        = 0x10006d2
	arabic_heh_goal         = 0x10006c1

	cyrillic_ghe_bar_upper        = 0x1000492
	cyrillic_ghe_bar              = 0x1000493
	cyrillic_zhe_descender_upper  = 0x1000496
	cyrillic_zhe_descender        = 0x1000497
	cyrillic_ka_descender_upper   = 0x100049a
	cyrillic_ka_descender         = 0x100049b
	cyrillic_ka_vertstroke_upper  = 0x100049c
	cyrillic_ka_vertstroke        = 0x100049d
	cyrillic_en_descender_upper   = 0x10004a2
	cyrillic_en_descender         = 0x10004a3
	cyrillic_u_straight_upper     = 0x10004ae
	cyrillic_u_straight           = 0x10004af
	cyrillic_u_straight_bar_upper = 0x10004b0
	cyrillic_u_straight_bar       = 0x10004b1
	cyrillic_ha_descender_upper   = 0x10004b2
	cyrillic_ha_descender         = 0x10004b3
	cyrillic_che_descender_upper  = 0x10004b6
	cyrillic_che_descender        = 0x10004b7
	cyrillic_che_vertstroke_upper = 0x10004b8
	cyrillic_che_vertstroke       = 0x10004b9
	cyrillic_shha_upper           = 0x10004ba
	cyrillic_shha                 = 0x10004bb

	cyrillic_schwa_upper    = 0x10004d8
	cyrillic_schwa          = 0x10004d9
	cyrillic_i_macron_upper = 0x10004e2
	cyrillic_i_macron       = 0x10004e3
	cyrillic_o_bar_upper    = 0x10004e8
	cyrillic_o_bar          = 0x10004e9
	cyrillic_u_macron_upper = 0x10004ee
	cyrillic_u_macron       = 0x10004ef

	serbian_dje                     = 0x06a1
	macedonia_gje                   = 0x06a2
	cyrillic_io                     = 0x06a3
	ukrainian_ie                    = 0x06a4
	macedonia_dse                   = 0x06a5
	ukrainian_i                     = 0x06a6
	ukrainian_yi                    = 0x06a7
	cyrillic_je                     = 0x06a8
	cyrillic_lje                    = 0x06a9
	cyrillic_nje                    = 0x06aa
	serbian_tshe                    = 0x06ab
	macedonia_kje                   = 0x06ac
	ukrainian_ghe_with_upturn       = 0x06ad
	byelorussian_shortu             = 0x06ae
	cyrillic_dzhe                   = 0x06af
	numerosign                      = 0x06b0
	serbian_dje_upper               = 0x06b1
	macedonia_gje_upper             = 0x06b2
	cyrillic_io_upper               = 0x06b3
	ukrainian_ie_upper              = 0x06b4
	macedonia_dse_upper             = 0x06b5
	ukrainian_i_upper               = 0x06b6
	ukrainian_yi_upper              = 0x06b7
	cyrillic_je_upper               = 0x06b8
	cyrillic_lje_upper              = 0x06b9
	cyrillic_nje_upper              = 0x06ba
	serbian_tshe_upper              = 0x06bb
	macedonia_kje_upper             = 0x06bc
	ukrainian_ghe_with_upturn_upper = 0x06bd
	byelorussian_shortu_upper       = 0x06be
	cyrillic_dzhe_upper             = 0x06bf
	cyrillic_yu                     = 0x06c0
	cyrillic_a                      = 0x06c1
	cyrillic_be                     = 0x06c2
	cyrillic_tse                    = 0x06c3
	cyrillic_de                     = 0x06c4
	cyrillic_ie                     = 0x06c5
	cyrillic_ef                     = 0x06c6
	cyrillic_ghe                    = 0x06c7
	cyrillic_ha                     = 0x06c8
	cyrillic_i                      = 0x06c9
	cyrillic_shorti                 = 0x06ca
	cyrillic_ka                     = 0x06cb
	cyrillic_el                     = 0x06cc
	cyrillic_em                     = 0x06cd
	cyrillic_en                     = 0x06ce
	cyrillic_o                      = 0x06cf
	cyrillic_pe                     = 0x06d0
	cyrillic_ya                     = 0x06d1
	cyrillic_er                     = 0x06d2
	cyrillic_es                     = 0x06d3
	cyrillic_te                     = 0x06d4
	cyrillic_u                      = 0x06d5
	cyrillic_zhe                    = 0x06d6
	cyrillic_ve                     = 0x06d7
	cyrillic_softsign               = 0x06d8
	cyrillic_yeru                   = 0x06d9
	cyrillic_ze                     = 0x06da
	cyrillic_sha                    = 0x06db
	cyrillic_e                      = 0x06dc
	cyrillic_shcha                  = 0x06dd
	cyrillic_che                    = 0x06de
	cyrillic_hardsign               = 0x06df
	cyrillic_yu_upper               = 0x06e0
	cyrillic_a_upper                = 0x06e1
	cyrillic_be_upper               = 0x06e2
	cyrillic_tse_upper              = 0x06e3
	cyrillic_de_upper               = 0x06e4
	cyrillic_ie_upper               = 0x06e5
	cyrillic_ef_upper               = 0x06e6
	cyrillic_ghe_upper              = 0x06e7
	cyrillic_ha_upper               = 0x06e8
	cyrillic_i_upper                = 0x06e9
	cyrillic_shorti_upper           = 0x06ea
	cyrillic_ka_upper               = 0x06eb
	cyrillic_el_upper               = 0x06ec
	cyrillic_em_upper               = 0x06ed
	cyrillic_en_upper               = 0x06ee
	cyrillic_o_upper                = 0x06ef
	cyrillic_pe_upper               = 0x06f0
	cyrillic_ya_upper               = 0x06f1
	cyrillic_er_upper               = 0x06f2
	cyrillic_es_upper               = 0x06f3
	cyrillic_te_upper               = 0x06f4
	cyrillic_u_upper                = 0x06f5
	cyrillic_zhe_upper              = 0x06f6
	cyrillic_ve_upper               = 0x06f7
	cyrillic_softsign_upper         = 0x06f8
	cyrillic_yeru_upper             = 0x06f9
	cyrillic_ze_upper               = 0x06fa
	cyrillic_sha_upper              = 0x06fb
	cyrillic_e_upper                = 0x06fc
	cyrillic_shcha_upper            = 0x06fd
	cyrillic_che_upper              = 0x06fe
	cyrillic_hardsign_upper         = 0x06ff
	greek_alphaaccent_upper         = 0x07a1
	greek_epsilonaccent_upper       = 0x07a2
	greek_etaaccent_upper           = 0x07a3
	greek_iotaaccent_upper          = 0x07a4
	greek_iotadieresis_upper        = 0x07a5
	greek_omicronaccent_upper       = 0x07a7
	greek_upsilonaccent_upper       = 0x07a8
	greek_upsilondieresis_upper     = 0x07a9
	greek_omegaaccent_upper         = 0x07ab
	greek_accentdieresis            = 0x07ae
	greek_horizbar                  = 0x07af
	greek_alphaaccent               = 0x07b1
	greek_epsilonaccent             = 0x07b2
	greek_etaaccent                 = 0x07b3
	greek_iotaaccent                = 0x07b4
	greek_iotadieresis              = 0x07b5
	greek_iotaaccentdieresis        = 0x07b6
	greek_omicronaccent             = 0x07b7
	greek_upsilonaccent             = 0x07b8
	greek_upsilondieresis           = 0x07b9
	greek_upsilonaccentdieresis     = 0x07ba
	greek_omegaaccent               = 0x07bb
	greek_alpha_upper               = 0x07c1
	greek_beta_upper                = 0x07c2
	greek_gamma_upper               = 0x07c3
	greek_delta_upper               = 0x07c4
	greek_epsilon_upper             = 0x07c5
	greek_zeta_upper                = 0x07c6
	greek_eta_upper                 = 0x07c7
	greek_theta_upper               = 0x07c8
	greek_iota_upper                = 0x07c9
	greek_kappa_upper               = 0x07ca
	greek_lamda_upper               = 0x07cb
	greek_mu_upper                  = 0x07cc
	greek_nu_upper                  = 0x07cd
	greek_xi_upper                  = 0x07ce
	greek_omicron_upper             = 0x07cf
	greek_pi_upper                  = 0x07d0
	greek_rho_upper                 = 0x07d1
	greek_sigma_upper               = 0x07d2
	greek_tau_upper                 = 0x07d4
	greek_upsilon_upper             = 0x07d5
	greek_phi_upper                 = 0x07d6
	greek_chi_upper                 = 0x07d7
	greek_psi_upper                 = 0x07d8
	greek_omega_upper               = 0x07d9
	greek_alpha                     = 0x07e1
	greek_beta                      = 0x07e2
	greek_gamma                     = 0x07e3
	greek_delta                     = 0x07e4
	greek_epsilon                   = 0x07e5
	greek_zeta                      = 0x07e6
	greek_eta                       = 0x07e7
	greek_theta                     = 0x07e8
	greek_iota                      = 0x07e9
	greek_kappa                     = 0x07ea
	greek_lamda                     = 0x07eb
	greek_mu                        = 0x07ec
	greek_nu                        = 0x07ed
	greek_xi                        = 0x07ee
	greek_omicron                   = 0x07ef
	greek_pi                        = 0x07f0
	greek_rho                       = 0x07f1
	greek_sigma                     = 0x07f2
	greek_finalsmallsigma           = 0x07f3
	greek_tau                       = 0x07f4
	greek_upsilon                   = 0x07f5
	greek_phi                       = 0x07f6
	greek_chi                       = 0x07f7
	greek_psi                       = 0x07f8
	greek_omega                     = 0x07f9
	leftradical                     = 0x08a1
	topleftradical                  = 0x08a2
	horizconnector                  = 0x08a3
	topintegral                     = 0x08a4
	botintegral                     = 0x08a5
	vertconnector                   = 0x08a6
	topleftsqbracket                = 0x08a7
	botleftsqbracket                = 0x08a8
	toprightsqbracket               = 0x08a9
	botrightsqbracket               = 0x08aa
	topleftparens                   = 0x08ab
	botleftparens                   = 0x08ac
	toprightparens                  = 0x08ad
	botrightparens                  = 0x08ae
	leftmiddlecurlybrace            = 0x08af
	rightmiddlecurlybrace           = 0x08b0
	topleftsummation                = 0x08b1
	botleftsummation                = 0x08b2
	topvertsummationconnector       = 0x08b3
	botvertsummationconnector       = 0x08b4
	toprightsummation               = 0x08b5
	botrightsummation               = 0x08b6
	rightmiddlesummation            = 0x08b7
	lessthanequal                   = 0x08bc
	notequal                        = 0x08bd
	greaterthanequal                = 0x08be
	integral                        = 0x08bf
	therefore                       = 0x08c0
	variation                       = 0x08c1
	infinity                        = 0x08c2
	nabla                           = 0x08c5
	approximate                     = 0x08c8
	similarequal                    = 0x08c9
	ifonlyif                        = 0x08cd
	implies                         = 0x08ce
	identical                       = 0x08cf
	radical                         = 0x08d6
	includedin                      = 0x08da
	includes                        = 0x08db
	intersection                    = 0x08dc
	union                           = 0x08dd
	logicaland                      = 0x08de
	logicalor                       = 0x08df
	partialderivative               = 0x08ef
	function                        = 0x08f6
	leftarrow                       = 0x08fb
	uparrow                         = 0x08fc
	rightarrow                      = 0x08fd
	downarrow                       = 0x08fe

	blank          = 0x09df
	soliddiamond   = 0x09e0
	checkerboard   = 0x09e1
	ht             = 0x09e2
	ff             = 0x09e3
	cr             = 0x09e4
	lf             = 0x09e5
	nl             = 0x09e8
	vt             = 0x09e9
	lowrightcorner = 0x09ea
	uprightcorner  = 0x09eb
	upleftcorner   = 0x09ec
	lowleftcorner  = 0x09ed
	crossinglines  = 0x09ee
	horizlinescan1 = 0x09ef
	horizlinescan3 = 0x09f0
	horizlinescan5 = 0x09f1
	horizlinescan7 = 0x09f2
	horizlinescan9 = 0x09f3
	leftt          = 0x09f4
	rightt         = 0x09f5
	bott           = 0x09f6
	topt           = 0x09f7
	vertbar        = 0x09f8

	emspace                = 0x0aa1
	enspace                = 0x0aa2
	em3space               = 0x0aa3
	em4space               = 0x0aa4
	digitspace             = 0x0aa5
	punctspace             = 0x0aa6
	thinspace              = 0x0aa7
	hairspace              = 0x0aa8
	emdash                 = 0x0aa9
	endash                 = 0x0aaa
	signifblank            = 0x0aac
	ellipsis               = 0x0aae
	doubbaselinedot        = 0x0aaf
	onethird               = 0x0ab0
	twothirds              = 0x0ab1
	onefifth               = 0x0ab2
	twofifths              = 0x0ab3
	threefifths            = 0x0ab4
	fourfifths             = 0x0ab5
	onesixth               = 0x0ab6
	fivesixths             = 0x0ab7
	careof                 = 0x0ab8
	figdash                = 0x0abb
	leftanglebracket       = 0x0abc
	decimalpoint           = 0x0abd
	rightanglebracket      = 0x0abe
	marker                 = 0x0abf
	oneeighth              = 0x0ac3
	threeeighths           = 0x0ac4
	fiveeighths            = 0x0ac5
	seveneighths           = 0x0ac6
	trademark              = 0x0ac9
	signaturemark          = 0x0aca
	trademarkincircle      = 0x0acb
	leftopentriangle       = 0x0acc
	rightopentriangle      = 0x0acd
	emopencircle           = 0x0ace
	emopenrectangle        = 0x0acf
	leftsinglequotemark    = 0x0ad0
	rightsinglequotemark   = 0x0ad1
	leftdoublequotemark    = 0x0ad2
	rightdoublequotemark   = 0x0ad3
	prescription           = 0x0ad4
	permille               = 0x0ad5
	minutes                = 0x0ad6
	seconds                = 0x0ad7
	latincross             = 0x0ad9
	hexagram               = 0x0ada
	filledrectbullet       = 0x0adb
	filledlefttribullet    = 0x0adc
	filledrighttribullet   = 0x0add
	emfilledcircle         = 0x0ade
	emfilledrect           = 0x0adf
	enopencircbullet       = 0x0ae0
	enopensquarebullet     = 0x0ae1
	openrectbullet         = 0x0ae2
	opentribulletup        = 0x0ae3
	opentribulletdown      = 0x0ae4
	openstar               = 0x0ae5
	enfilledcircbullet     = 0x0ae6
	enfilledsqbullet       = 0x0ae7
	filledtribulletup      = 0x0ae8
	filledtribulletdown    = 0x0ae9
	leftpointer            = 0x0aea
	rightpointer           = 0x0aeb
	club                   = 0x0aec
	diamond                = 0x0aed
	heart                  = 0x0aee
	maltesecross           = 0x0af0
	dagger                 = 0x0af1
	doubledagger           = 0x0af2
	checkmark              = 0x0af3
	ballotcross            = 0x0af4
	musicalsharp           = 0x0af5
	musicalflat            = 0x0af6
	malesymbol             = 0x0af7
	femalesymbol           = 0x0af8
	telephone              = 0x0af9
	telephonerecorder      = 0x0afa
	phonographcopyright    = 0x0afb
	caret                  = 0x0afc
	singlelowquotemark     = 0x0afd
	doublelowquotemark     = 0x0afe
	cursor                 = 0x0aff
	leftcaret              = 0x0ba3
	rightcaret             = 0x0ba6
	downcaret              = 0x0ba8
	upcaret                = 0x0ba9
	overbar                = 0x0bc0
	downtack               = 0x0bc2
	upshoe                 = 0x0bc3
	downstile              = 0x0bc4
	underbar               = 0x0bc6
	jot                    = 0x0bca
	quad                   = 0x0bcc
	uptack                 = 0x0bce
	circle                 = 0x0bcf
	upstile                = 0x0bd3
	downshoe               = 0x0bd6
	rightshoe              = 0x0bd8
	leftshoe               = 0x0bda
	lefttack               = 0x0bdc
	righttack              = 0x0bfc
	hebrew_doublelowline   = 0x0cdf
	hebrew_aleph           = 0x0ce0
	hebrew_bet             = 0x0ce1
	hebrew_gimel           = 0x0ce2
	hebrew_dalet           = 0x0ce3
	hebrew_he              = 0x0ce4
	hebrew_waw             = 0x0ce5
	hebrew_zain            = 0x0ce6
	hebrew_chet            = 0x0ce7
	hebrew_tet             = 0x0ce8
	hebrew_yod             = 0x0ce9
	hebrew_finalkaph       = 0x0cea
	hebrew_kaph            = 0x0ceb
	hebrew_lamed           = 0x0cec
	hebrew_finalmem        = 0x0ced
	hebrew_mem             = 0x0cee
	hebrew_finalnun        = 0x0cef
	hebrew_nun             = 0x0cf0
	hebrew_samech          = 0x0cf1
	hebrew_ayin            = 0x0cf2
	hebrew_finalpe         = 0x0cf3
	hebrew_pe              = 0x0cf4
	hebrew_finalzade       = 0x0cf5
	hebrew_zade            = 0x0cf6
	hebrew_qoph            = 0x0cf7
	hebrew_resh            = 0x0cf8
	hebrew_shin            = 0x0cf9
	hebrew_taw             = 0x0cfa
	thai_kokai             = 0x0da1
	thai_khokhai           = 0x0da2
	thai_khokhuat          = 0x0da3
	thai_khokhwai          = 0x0da4
	thai_khokhon           = 0x0da5
	thai_khorakhang        = 0x0da6
	thai_ngongu            = 0x0da7
	thai_chochan           = 0x0da8
	thai_choching          = 0x0da9
	thai_chochang          = 0x0daa
	thai_soso              = 0x0dab
	thai_chochoe           = 0x0dac
	thai_yoying            = 0x0dad
	thai_dochada           = 0x0dae
	thai_topatak           = 0x0daf
	thai_thothan           = 0x0db0
	thai_thonangmontho     = 0x0db1
	thai_thophuthao        = 0x0db2
	thai_nonen             = 0x0db3
	thai_dodek             = 0x0db4
	thai_totao             = 0x0db5
	thai_thothung          = 0x0db6
	thai_thothahan         = 0x0db7
	thai_thothong          = 0x0db8
	thai_nonu              = 0x0db9
	thai_bobaimai          = 0x0dba
	thai_popla             = 0x0dbb
	thai_phophung          = 0x0dbc
	thai_fofa              = 0x0dbd
	thai_phophan           = 0x0dbe
	thai_fofan             = 0x0dbf
	thai_phosamphao        = 0x0dc0
	thai_moma              = 0x0dc1
	thai_yoyak             = 0x0dc2
	thai_rorua             = 0x0dc3
	thai_ru                = 0x0dc4
	thai_loling            = 0x0dc5
	thai_lu                = 0x0dc6
	thai_wowaen            = 0x0dc7
	thai_sosala            = 0x0dc8
	thai_sorusi            = 0x0dc9
	thai_sosua             = 0x0dca
	thai_hohip             = 0x0dcb
	thai_lochula           = 0x0dcc
	thai_oang              = 0x0dcd
	thai_honokhuk          = 0x0dce
	thai_paiyannoi         = 0x0dcf
	thai_saraa             = 0x0dd0
	thai_maihanakat        = 0x0dd1
	thai_saraaa            = 0x0dd2
	thai_saraam            = 0x0dd3
	thai_sarai             = 0x0dd4
	thai_saraii            = 0x0dd5
	thai_saraue            = 0x0dd6
	thai_sarauee           = 0x0dd7
	thai_sarau             = 0x0dd8
	thai_sarauu            = 0x0dd9
	thai_phinthu           = 0x0dda
	thai_maihanakat_maitho = 0x0dde
	thai_baht              = 0x0ddf
	thai_sarae             = 0x0de0
	thai_saraae            = 0x0de1
	thai_sarao             = 0x0de2
	thai_saraaimaimuan     = 0x0de3
	thai_saraaimaimalai    = 0x0de4
	thai_lakkhangyao       = 0x0de5
	thai_maiyamok          = 0x0de6
	thai_maitaikhu         = 0x0de7
	thai_maiek             = 0x0de8
	thai_maitho            = 0x0de9
	thai_maitri            = 0x0dea
	thai_maichattawa       = 0x0deb
	thai_thanthakhat       = 0x0dec
	thai_nikhahit          = 0x0ded
	thai_leksun            = 0x0df0
	thai_leknung           = 0x0df1
	thai_leksong           = 0x0df2
	thai_leksam            = 0x0df3
	thai_leksi             = 0x0df4
	thai_lekha             = 0x0df5
	thai_lekhok            = 0x0df6
	thai_lekchet           = 0x0df7
	thai_lekpaet           = 0x0df8
	thai_lekkao            = 0x0df9

	hangul           = 0xff31
	hangul_start     = 0xff32
	hangul_end       = 0xff33
	hangul_hanja     = 0xff34
	hangul_jamo      = 0xff35
	hangul_romaja    = 0xff36
	hangul_jeonja    = 0xff38
	hangul_banja     = 0xff39
	hangul_prehanja  = 0xff3a
	hangul_posthanja = 0xff3b
	hangul_special   = 0xff3f

	hangul_kiyeog      = 0x0ea1
	hangul_ssangkiyeog = 0x0ea2
	hangul_kiyeogsios  = 0x0ea3
	hangul_nieun       = 0x0ea4
	hangul_nieunjieuj  = 0x0ea5
	hangul_nieunhieuh  = 0x0ea6
	hangul_dikeud      = 0x0ea7
	hangul_ssangdikeud = 0x0ea8
	hangul_rieul       = 0x0ea9
	hangul_rieulkiyeog = 0x0eaa
	hangul_rieulmieum  = 0x0eab
	hangul_rieulpieub  = 0x0eac
	hangul_rieulsios   = 0x0ead
	hangul_rieultieut  = 0x0eae
	hangul_rieulphieuf = 0x0eaf
	hangul_rieulhieuh  = 0x0eb0
	hangul_mieum       = 0x0eb1
	hangul_pieub       = 0x0eb2
	hangul_ssangpieub  = 0x0eb3
	hangul_pieubsios   = 0x0eb4
	hangul_sios        = 0x0eb5
	hangul_ssangsios   = 0x0eb6
	hangul_ieung       = 0x0eb7
	hangul_jieuj       = 0x0eb8
	hangul_ssangjieuj  = 0x0eb9
	hangul_cieuc       = 0x0eba
	hangul_khieuq      = 0x0ebb
	hangul_tieut       = 0x0ebc
	hangul_phieuf      = 0x0ebd
	hangul_hieuh       = 0x0ebe

	hangul_a   = 0x0ebf
	hangul_ae  = 0x0ec0
	hangul_ya  = 0x0ec1
	hangul_yae = 0x0ec2
	hangul_eo  = 0x0ec3
	hangul_e   = 0x0ec4
	hangul_yeo = 0x0ec5
	hangul_ye  = 0x0ec6
	hangul_o   = 0x0ec7
	hangul_wa  = 0x0ec8
	hangul_wae = 0x0ec9
	hangul_oe  = 0x0eca
	hangul_yo  = 0x0ecb
	hangul_u   = 0x0ecc
	hangul_weo = 0x0ecd
	hangul_we  = 0x0ece
	hangul_wi  = 0x0ecf
	hangul_yu  = 0x0ed0
	hangul_eu  = 0x0ed1
	hangul_yi  = 0x0ed2
	hangul_i   = 0x0ed3

	hangul_j_kiyeog      = 0x0ed4
	hangul_j_ssangkiyeog = 0x0ed5
	hangul_j_kiyeogsios  = 0x0ed6
	hangul_j_nieun       = 0x0ed7
	hangul_j_nieunjieuj  = 0x0ed8
	hangul_j_nieunhieuh  = 0x0ed9
	hangul_j_dikeud      = 0x0eda
	hangul_j_rieul       = 0x0edb
	hangul_j_rieulkiyeog = 0x0edc
	hangul_j_rieulmieum  = 0x0edd
	hangul_j_rieulpieub  = 0x0ede
	hangul_j_rieulsios   = 0x0edf
	hangul_j_rieultieut  = 0x0ee0
	hangul_j_rieulphieuf = 0x0ee1
	hangul_j_rieulhieuh  = 0x0ee2
	hangul_j_mieum       = 0x0ee3
	hangul_j_pieub       = 0x0ee4
	hangul_j_pieubsios   = 0x0ee5
	hangul_j_sios        = 0x0ee6
	hangul_j_ssangsios   = 0x0ee7
	hangul_j_ieung       = 0x0ee8
	hangul_j_jieuj       = 0x0ee9
	hangul_j_cieuc       = 0x0eea
	hangul_j_khieuq      = 0x0eeb
	hangul_j_tieut       = 0x0eec
	hangul_j_phieuf      = 0x0eed
	hangul_j_hieuh       = 0x0eee

	hangul_rieulyeorinhieuh   = 0x0eef
	hangul_sunkyeongeummieum  = 0x0ef0
	hangul_sunkyeongeumpieub  = 0x0ef1
	hangul_pansios            = 0x0ef2
	hangul_kkogjidalrinieung  = 0x0ef3
	hangul_sunkyeongeumphieuf = 0x0ef4
	hangul_yeorinhieuh        = 0x0ef5

	hangul_araea  = 0x0ef6
	hangul_araeae = 0x0ef7

	hangul_j_pansios           = 0x0ef8
	hangul_j_kkogjidalrinieung = 0x0ef9
	hangul_j_yeorinhieuh       = 0x0efa

	korean_won = 0x0eff

	armenian_ligature_ew     = 0x1000587
	armenian_full_stop       = 0x1000589
	armenian_separation_mark = 0x100055d
	armenian_hyphen          = 0x100058a
	armenian_exclam          = 0x100055c
	armenian_accent          = 0x100055b
	armenian_question        = 0x100055e
	armenian_ayb_upper       = 0x1000531
	armenian_ayb             = 0x1000561
	armenian_ben_upper       = 0x1000532
	armenian_ben             = 0x1000562
	armenian_gim_upper       = 0x1000533
	armenian_gim             = 0x1000563
	armenian_da_upper        = 0x1000534
	armenian_da              = 0x1000564
	armenian_yech_upper      = 0x1000535
	armenian_yech            = 0x1000565
	armenian_za_upper        = 0x1000536
	armenian_za              = 0x1000566
	armenian_e_upper         = 0x1000537
	armenian_e               = 0x1000567
	armenian_at_upper        = 0x1000538
	armenian_at              = 0x1000568
	armenian_to_upper        = 0x1000539
	armenian_to              = 0x1000569
	armenian_zhe_upper       = 0x100053a
	armenian_zhe             = 0x100056a
	armenian_ini_upper       = 0x100053b
	armenian_ini             = 0x100056b
	armenian_lyun_upper      = 0x100053c
	armenian_lyun            = 0x100056c
	armenian_khe_upper       = 0x100053d
	armenian_khe             = 0x100056d
	armenian_tsa_upper       = 0x100053e
	armenian_tsa             = 0x100056e
	armenian_ken_upper       = 0x100053f
	armenian_ken             = 0x100056f
	armenian_ho_upper        = 0x1000540
	armenian_ho              = 0x1000570
	armenian_dza_upper       = 0x1000541
	armenian_dza             = 0x1000571
	armenian_ghat_upper      = 0x1000542
	armenian_ghat            = 0x1000572
	armenian_tche_upper      = 0x1000543
	armenian_tche            = 0x1000573
	armenian_men_upper       = 0x1000544
	armenian_men             = 0x1000574
	armenian_hi_upper        = 0x1000545
	armenian_hi              = 0x1000575
	armenian_nu_upper        = 0x1000546
	armenian_nu              = 0x1000576
	armenian_sha_upper       = 0x1000547
	armenian_sha             = 0x1000577
	armenian_vo_upper        = 0x1000548
	armenian_vo              = 0x1000578
	armenian_cha_upper       = 0x1000549
	armenian_cha             = 0x1000579
	armenian_pe_upper        = 0x100054a
	armenian_pe              = 0x100057a
	armenian_je_upper        = 0x100054b
	armenian_je              = 0x100057b
	armenian_ra_upper        = 0x100054c
	armenian_ra              = 0x100057c
	armenian_se_upper        = 0x100054d
	armenian_se              = 0x100057d
	armenian_vev_upper       = 0x100054e
	armenian_vev             = 0x100057e
	armenian_tyun_upper      = 0x100054f
	armenian_tyun            = 0x100057f
	armenian_re_upper        = 0x1000550
	armenian_re              = 0x1000580
	armenian_tso_upper       = 0x1000551
	armenian_tso             = 0x1000581
	armenian_vyun_upper      = 0x1000552
	armenian_vyun            = 0x1000582
	armenian_pyur_upper      = 0x1000553
	armenian_pyur            = 0x1000583
	armenian_ke_upper        = 0x1000554
	armenian_ke              = 0x1000584
	armenian_o_upper         = 0x1000555
	armenian_o               = 0x1000585
	armenian_fe_upper        = 0x1000556
	armenian_fe              = 0x1000586
	armenian_apostrophe      = 0x100055a
	georgian_an              = 0x10010d0
	georgian_ban             = 0x10010d1
	georgian_gan             = 0x10010d2
	georgian_don             = 0x10010d3
	georgian_en              = 0x10010d4
	georgian_vin             = 0x10010d5
	georgian_zen             = 0x10010d6
	georgian_tan             = 0x10010d7
	georgian_in              = 0x10010d8
	georgian_kan             = 0x10010d9
	georgian_las             = 0x10010da
	georgian_man             = 0x10010db
	georgian_nar             = 0x10010dc
	georgian_on              = 0x10010dd
	georgian_par             = 0x10010de
	georgian_zhar            = 0x10010df
	georgian_rae             = 0x10010e0
	georgian_san             = 0x10010e1
	georgian_tar             = 0x10010e2
	georgian_un              = 0x10010e3
	georgian_phar            = 0x10010e4
	georgian_khar            = 0x10010e5
	georgian_ghan            = 0x10010e6
	georgian_qar             = 0x10010e7
	georgian_shin            = 0x10010e8
	georgian_chin            = 0x10010e9
	georgian_can             = 0x10010ea
	georgian_jil             = 0x10010eb
	georgian_cil             = 0x10010ec
	georgian_char            = 0x10010ed
	georgian_xan             = 0x10010ee
	georgian_jhan            = 0x10010ef
	georgian_hae             = 0x10010f0
	georgian_he              = 0x10010f1
	georgian_hie             = 0x10010f2
	georgian_we              = 0x10010f3
	georgian_har             = 0x10010f4
	georgian_hoe             = 0x10010f5
	georgian_fi              = 0x10010f6

	xabovedot_upper = 0x1001e8a
	ibreve_upper    = 0x100012c
	zstroke_upper   = 0x10001b5
	gcaron_upper    = 0x10001e6
	ocaron_upper    = 0x10001d1
	obarred_upper   = 0x100019f
	xabovedot       = 0x1001e8b
	ibreve          = 0x100012d
	zstroke         = 0x10001b6
	gcaron          = 0x10001e7
	ocaron          = 0x10001d2
	obarred         = 0x1000275
	schwa_upper     = 0x100018f
	schwa           = 0x1000259
	ezh_upper       = 0x10001b7
	ezh             = 0x1000292

	lbelowdot_upper = 0x1001e36
	lbelowdot       = 0x1001e37

	abelowdot_upper           = 0x1001ea0
	abelowdot                 = 0x1001ea1
	ahook_upper               = 0x1001ea2
	ahook                     = 0x1001ea3
	acircumflexacute_upper    = 0x1001ea4
	acircumflexacute          = 0x1001ea5
	acircumflexgrave_upper    = 0x1001ea6
	acircumflexgrave          = 0x1001ea7
	acircumflexhook_upper     = 0x1001ea8
	acircumflexhook           = 0x1001ea9
	acircumflextilde_upper    = 0x1001eaa
	acircumflextilde          = 0x1001eab
	acircumflexbelowdot_upper = 0x1001eac
	acircumflexbelowdot       = 0x1001ead
	abreveacute_upper         = 0x1001eae
	abreveacute               = 0x1001eaf
	abrevegrave_upper         = 0x1001eb0
	abrevegrave               = 0x1001eb1
	abrevehook_upper          = 0x1001eb2
	abrevehook                = 0x1001eb3
	abrevetilde_upper         = 0x1001eb4
	abrevetilde               = 0x1001eb5
	abrevebelowdot_upper      = 0x1001eb6
	abrevebelowdot            = 0x1001eb7
	ebelowdot_upper           = 0x1001eb8
	ebelowdot                 = 0x1001eb9
	ehook_upper               = 0x1001eba
	ehook                     = 0x1001ebb
	etilde_upper              = 0x1001ebc
	etilde                    = 0x1001ebd
	ecircumflexacute_upper    = 0x1001ebe
	ecircumflexacute          = 0x1001ebf
	ecircumflexgrave_upper    = 0x1001ec0
	ecircumflexgrave          = 0x1001ec1
	ecircumflexhook_upper     = 0x1001ec2
	ecircumflexhook           = 0x1001ec3
	ecircumflextilde_upper    = 0x1001ec4
	ecircumflextilde          = 0x1001ec5
	ecircumflexbelowdot_upper = 0x1001ec6
	ecircumflexbelowdot       = 0x1001ec7
	ihook_upper               = 0x1001ec8
	ihook                     = 0x1001ec9
	ibelowdot_upper           = 0x1001eca
	ibelowdot                 = 0x1001ecb
	obelowdot_upper           = 0x1001ecc
	obelowdot                 = 0x1001ecd
	ohook_upper               = 0x1001ece
	ohook                     = 0x1001ecf
	ocircumflexacute_upper    = 0x1001ed0
	ocircumflexacute          = 0x1001ed1
	ocircumflexgrave_upper    = 0x1001ed2
	ocircumflexgrave          = 0x1001ed3
	ocircumflexhook_upper     = 0x1001ed4
	ocircumflexhook           = 0x1001ed5
	ocircumflextilde_upper    = 0x1001ed6
	ocircumflextilde          = 0x1001ed7
	ocircumflexbelowdot_upper = 0x1001ed8
	ocircumflexbelowdot       = 0x1001ed9
	ohornacute_upper          = 0x1001eda
	ohornacute                = 0x1001edb
	ohorngrave_upper          = 0x1001edc
	ohorngrave                = 0x1001edd
	ohornhook_upper           = 0x1001ede
	ohornhook                 = 0x1001edf
	ohorntilde_upper          = 0x1001ee0
	ohorntilde                = 0x1001ee1
	ohornbelowdot_upper       = 0x1001ee2
	ohornbelowdot             = 0x1001ee3
	ubelowdot_upper           = 0x1001ee4
	ubelowdot                 = 0x1001ee5
	uhook_upper               = 0x1001ee6
	uhook                     = 0x1001ee7
	uhornacute_upper          = 0x1001ee8
	uhornacute                = 0x1001ee9
	uhorngrave_upper          = 0x1001eea
	uhorngrave                = 0x1001eeb
	uhornhook_upper           = 0x1001eec
	uhornhook                 = 0x1001eed
	uhorntilde_upper          = 0x1001eee
	uhorntilde                = 0x1001eef
	uhornbelowdot_upper       = 0x1001ef0
	uhornbelowdot             = 0x1001ef1
	ybelowdot_upper           = 0x1001ef4
	ybelowdot                 = 0x1001ef5
	yhook_upper               = 0x1001ef6
	yhook                     = 0x1001ef7
	ytilde_upper              = 0x1001ef8
	ytilde                    = 0x1001ef9
	ohorn_upper               = 0x10001a0
	ohorn                     = 0x10001a1
	uhorn_upper               = 0x10001af
	uhorn                     = 0x10001b0
	combining_tilde           = 0x1000303
	combining_grave           = 0x1000300
	combining_acute           = 0x1000301
	combining_hook            = 0x1000309
	combining_belowdot        = 0x1000323

	ecusign       = 0x10020a0
	colonsign     = 0x10020a1
	cruzeirosign  = 0x10020a2
	ffrancsign    = 0x10020a3
	lirasign      = 0x10020a4
	millsign      = 0x10020a5
	nairasign     = 0x10020a6
	pesetasign    = 0x10020a7
	rupeesign     = 0x10020a8
	wonsign       = 0x10020a9
	newsheqelsign = 0x10020aa
	dongsign      = 0x10020ab
	eurosign      = 0x20ac

	zerosuperior     = 0x1002070
	foursuperior     = 0x1002074
	fivesuperior     = 0x1002075
	sixsuperior      = 0x1002076
	sevensuperior    = 0x1002077
	eightsuperior    = 0x1002078
	ninesuperior     = 0x1002079
	zerosubscript    = 0x1002080
	onesubscript     = 0x1002081
	twosubscript     = 0x1002082
	threesubscript   = 0x1002083
	foursubscript    = 0x1002084
	fivesubscript    = 0x1002085
	sixsubscript     = 0x1002086
	sevensubscript   = 0x1002087
	eightsubscript   = 0x1002088
	ninesubscript    = 0x1002089
	partdifferential = 0x1002202
	emptyset         = 0x1002205
	elementof        = 0x1002208
	notelementof     = 0x1002209
	containsas       = 0x100220b
	squareroot       = 0x100221a
	cuberoot         = 0x100221b
	fourthroot       = 0x100221c
	dintegral        = 0x100222c
	tintegral        = 0x100222d
	because          = 0x1002235
	approxeq         = 0x1002248
	notapproxeq      = 0x1002247
	notidentical     = 0x1002262
	stricteq         = 0x1002263

	braille_dot_1         = 0xfff1
	braille_dot_2         = 0xfff2
	braille_dot_3         = 0xfff3
	braille_dot_4         = 0xfff4
	braille_dot_5         = 0xfff5
	braille_dot_6         = 0xfff6
	braille_dot_7         = 0xfff7
	braille_dot_8         = 0xfff8
	braille_dot_9         = 0xfff9
	braille_dot_10        = 0xfffa
	braille_blank         = 0x1002800
	braille_dots_1        = 0x1002801
	braille_dots_2        = 0x1002802
	braille_dots_12       = 0x1002803
	braille_dots_3        = 0x1002804
	braille_dots_13       = 0x1002805
	braille_dots_23       = 0x1002806
	braille_dots_123      = 0x1002807
	braille_dots_4        = 0x1002808
	braille_dots_14       = 0x1002809
	braille_dots_24       = 0x100280a
	braille_dots_124      = 0x100280b
	braille_dots_34       = 0x100280c
	braille_dots_134      = 0x100280d
	braille_dots_234      = 0x100280e
	braille_dots_1234     = 0x100280f
	braille_dots_5        = 0x1002810
	braille_dots_15       = 0x1002811
	braille_dots_25       = 0x1002812
	braille_dots_125      = 0x1002813
	braille_dots_35       = 0x1002814
	braille_dots_135      = 0x1002815
	braille_dots_235      = 0x1002816
	braille_dots_1235     = 0x1002817
	braille_dots_45       = 0x1002818
	braille_dots_145      = 0x1002819
	braille_dots_245      = 0x100281a
	braille_dots_1245     = 0x100281b
	braille_dots_345      = 0x100281c
	braille_dots_1345     = 0x100281d
	braille_dots_2345     = 0x100281e
	braille_dots_12345    = 0x100281f
	braille_dots_6        = 0x1002820
	braille_dots_16       = 0x1002821
	braille_dots_26       = 0x1002822
	braille_dots_126      = 0x1002823
	braille_dots_36       = 0x1002824
	braille_dots_136      = 0x1002825
	braille_dots_236      = 0x1002826
	braille_dots_1236     = 0x1002827
	braille_dots_46       = 0x1002828
	braille_dots_146      = 0x1002829
	braille_dots_246      = 0x100282a
	braille_dots_1246     = 0x100282b
	braille_dots_346      = 0x100282c
	braille_dots_1346     = 0x100282d
	braille_dots_2346     = 0x100282e
	braille_dots_12346    = 0x100282f
	braille_dots_56       = 0x1002830
	braille_dots_156      = 0x1002831
	braille_dots_256      = 0x1002832
	braille_dots_1256     = 0x1002833
	braille_dots_356      = 0x1002834
	braille_dots_1356     = 0x1002835
	braille_dots_2356     = 0x1002836
	braille_dots_12356    = 0x1002837
	braille_dots_456      = 0x1002838
	braille_dots_1456     = 0x1002839
	braille_dots_2456     = 0x100283a
	braille_dots_12456    = 0x100283b
	braille_dots_3456     = 0x100283c
	braille_dots_13456    = 0x100283d
	braille_dots_23456    = 0x100283e
	braille_dots_123456   = 0x100283f
	braille_dots_7        = 0x1002840
	braille_dots_17       = 0x1002841
	braille_dots_27       = 0x1002842
	braille_dots_127      = 0x1002843
	braille_dots_37       = 0x1002844
	braille_dots_137      = 0x1002845
	braille_dots_237      = 0x1002846
	braille_dots_1237     = 0x1002847
	braille_dots_47       = 0x1002848
	braille_dots_147      = 0x1002849
	braille_dots_247      = 0x100284a
	braille_dots_1247     = 0x100284b
	braille_dots_347      = 0x100284c
	braille_dots_1347     = 0x100284d
	braille_dots_2347     = 0x100284e
	braille_dots_12347    = 0x100284f
	braille_dots_57       = 0x1002850
	braille_dots_157      = 0x1002851
	braille_dots_257      = 0x1002852
	braille_dots_1257     = 0x1002853
	braille_dots_357      = 0x1002854
	braille_dots_1357     = 0x1002855
	braille_dots_2357     = 0x1002856
	braille_dots_12357    = 0x1002857
	braille_dots_457      = 0x1002858
	braille_dots_1457     = 0x1002859
	braille_dots_2457     = 0x100285a
	braille_dots_12457    = 0x100285b
	braille_dots_3457     = 0x100285c
	braille_dots_13457    = 0x100285d
	braille_dots_23457    = 0x100285e
	braille_dots_123457   = 0x100285f
	braille_dots_67       = 0x1002860
	braille_dots_167      = 0x1002861
	braille_dots_267      = 0x1002862
	braille_dots_1267     = 0x1002863
	braille_dots_367      = 0x1002864
	braille_dots_1367     = 0x1002865
	braille_dots_2367     = 0x1002866
	braille_dots_12367    = 0x1002867
	braille_dots_467      = 0x1002868
	braille_dots_1467     = 0x1002869
	braille_dots_2467     = 0x100286a
	braille_dots_12467    = 0x100286b
	braille_dots_3467     = 0x100286c
	braille_dots_13467    = 0x100286d
	braille_dots_23467    = 0x100286e
	braille_dots_123467   = 0x100286f
	braille_dots_567      = 0x1002870
	braille_dots_1567     = 0x1002871
	braille_dots_2567     = 0x1002872
	braille_dots_12567    = 0x1002873
	braille_dots_3567     = 0x1002874
	braille_dots_13567    = 0x1002875
	braille_dots_23567    = 0x1002876
	braille_dots_123567   = 0x1002877
	braille_dots_4567     = 0x1002878
	braille_dots_14567    = 0x1002879
	braille_dots_24567    = 0x100287a
	braille_dots_124567   = 0x100287b
	braille_dots_34567    = 0x100287c
	braille_dots_134567   = 0x100287d
	braille_dots_234567   = 0x100287e
	braille_dots_1234567  = 0x100287f
	braille_dots_8        = 0x1002880
	braille_dots_18       = 0x1002881
	braille_dots_28       = 0x1002882
	braille_dots_128      = 0x1002883
	braille_dots_38       = 0x1002884
	braille_dots_138      = 0x1002885
	braille_dots_238      = 0x1002886
	braille_dots_1238     = 0x1002887
	braille_dots_48       = 0x1002888
	braille_dots_148      = 0x1002889
	braille_dots_248      = 0x100288a
	braille_dots_1248     = 0x100288b
	braille_dots_348      = 0x100288c
	braille_dots_1348     = 0x100288d
	braille_dots_2348     = 0x100288e
	braille_dots_12348    = 0x100288f
	braille_dots_58       = 0x1002890
	braille_dots_158      = 0x1002891
	braille_dots_258      = 0x1002892
	braille_dots_1258     = 0x1002893
	braille_dots_358      = 0x1002894
	braille_dots_1358     = 0x1002895
	braille_dots_2358     = 0x1002896
	braille_dots_12358    = 0x1002897
	braille_dots_458      = 0x1002898
	braille_dots_1458     = 0x1002899
	braille_dots_2458     = 0x100289a
	braille_dots_12458    = 0x100289b
	braille_dots_3458     = 0x100289c
	braille_dots_13458    = 0x100289d
	braille_dots_23458    = 0x100289e
	braille_dots_123458   = 0x100289f
	braille_dots_68       = 0x10028a0
	braille_dots_168      = 0x10028a1
	braille_dots_268      = 0x10028a2
	braille_dots_1268     = 0x10028a3
	braille_dots_368      = 0x10028a4
	braille_dots_1368     = 0x10028a5
	braille_dots_2368     = 0x10028a6
	braille_dots_12368    = 0x10028a7
	braille_dots_468      = 0x10028a8
	braille_dots_1468     = 0x10028a9
	braille_dots_2468     = 0x10028aa
	braille_dots_12468    = 0x10028ab
	braille_dots_3468     = 0x10028ac
	braille_dots_13468    = 0x10028ad
	braille_dots_23468    = 0x10028ae
	braille_dots_123468   = 0x10028af
	braille_dots_568      = 0x10028b0
	braille_dots_1568     = 0x10028b1
	braille_dots_2568     = 0x10028b2
	braille_dots_12568    = 0x10028b3
	braille_dots_3568     = 0x10028b4
	braille_dots_13568    = 0x10028b5
	braille_dots_23568    = 0x10028b6
	braille_dots_123568   = 0x10028b7
	braille_dots_4568     = 0x10028b8
	braille_dots_14568    = 0x10028b9
	braille_dots_24568    = 0x10028ba
	braille_dots_124568   = 0x10028bb
	braille_dots_34568    = 0x10028bc
	braille_dots_134568   = 0x10028bd
	braille_dots_234568   = 0x10028be
	braille_dots_1234568  = 0x10028bf
	braille_dots_78       = 0x10028c0
	braille_dots_178      = 0x10028c1
	braille_dots_278      = 0x10028c2
	braille_dots_1278     = 0x10028c3
	braille_dots_378      = 0x10028c4
	braille_dots_1378     = 0x10028c5
	braille_dots_2378     = 0x10028c6
	braille_dots_12378    = 0x10028c7
	braille_dots_478      = 0x10028c8
	braille_dots_1478     = 0x10028c9
	braille_dots_2478     = 0x10028ca
	braille_dots_12478    = 0x10028cb
	braille_dots_3478     = 0x10028cc
	braille_dots_13478    = 0x10028cd
	braille_dots_23478    = 0x10028ce
	braille_dots_123478   = 0x10028cf
	braille_dots_578      = 0x10028d0
	braille_dots_1578     = 0x10028d1
	braille_dots_2578     = 0x10028d2
	braille_dots_12578    = 0x10028d3
	braille_dots_3578     = 0x10028d4
	braille_dots_13578    = 0x10028d5
	braille_dots_23578    = 0x10028d6
	braille_dots_123578   = 0x10028d7
	braille_dots_4578     = 0x10028d8
	braille_dots_14578    = 0x10028d9
	braille_dots_24578    = 0x10028da
	braille_dots_124578   = 0x10028db
	braille_dots_34578    = 0x10028dc
	braille_dots_134578   = 0x10028dd
	braille_dots_234578   = 0x10028de
	braille_dots_1234578  = 0x10028df
	braille_dots_678      = 0x10028e0
	braille_dots_1678     = 0x10028e1
	braille_dots_2678     = 0x10028e2
	braille_dots_12678    = 0x10028e3
	braille_dots_3678     = 0x10028e4
	braille_dots_13678    = 0x10028e5
	braille_dots_23678    = 0x10028e6
	braille_dots_123678   = 0x10028e7
	braille_dots_4678     = 0x10028e8
	braille_dots_14678    = 0x10028e9
	braille_dots_24678    = 0x10028ea
	braille_dots_124678   = 0x10028eb
	braille_dots_34678    = 0x10028ec
	braille_dots_134678   = 0x10028ed
	braille_dots_234678   = 0x10028ee
	braille_dots_1234678  = 0x10028ef
	braille_dots_5678     = 0x10028f0
	braille_dots_15678    = 0x10028f1
	braille_dots_25678    = 0x10028f2
	braille_dots_125678   = 0x10028f3
	braille_dots_35678    = 0x10028f4
	braille_dots_135678   = 0x10028f5
	braille_dots_235678   = 0x10028f6
	braille_dots_1235678  = 0x10028f7
	braille_dots_45678    = 0x10028f8
	braille_dots_145678   = 0x10028f9
	braille_dots_245678   = 0x10028fa
	braille_dots_1245678  = 0x10028fb
	braille_dots_345678   = 0x10028fc
	braille_dots_1345678  = 0x10028fd
	braille_dots_2345678  = 0x10028fe
	braille_dots_12345678 = 0x10028ff

	sinh_ng         = 0x1000d82
	sinh_h2         = 0x1000d83
	sinh_a          = 0x1000d85
	sinh_aa         = 0x1000d86
	sinh_ae         = 0x1000d87
	sinh_aee        = 0x1000d88
	sinh_i          = 0x1000d89
	sinh_ii         = 0x1000d8a
	sinh_u          = 0x1000d8b
	sinh_uu         = 0x1000d8c
	sinh_ri         = 0x1000d8d
	sinh_rii        = 0x1000d8e
	sinh_lu         = 0x1000d8f
	sinh_luu        = 0x1000d90
	sinh_e          = 0x1000d91
	sinh_ee         = 0x1000d92
	sinh_ai         = 0x1000d93
	sinh_o          = 0x1000d94
	sinh_oo         = 0x1000d95
	sinh_au         = 0x1000d96
	sinh_ka         = 0x1000d9a
	sinh_kha        = 0x1000d9b
	sinh_ga         = 0x1000d9c
	sinh_gha        = 0x1000d9d
	sinh_ng2        = 0x1000d9e
	sinh_nga        = 0x1000d9f
	sinh_ca         = 0x1000da0
	sinh_cha        = 0x1000da1
	sinh_ja         = 0x1000da2
	sinh_jha        = 0x1000da3
	sinh_nya        = 0x1000da4
	sinh_jnya       = 0x1000da5
	sinh_nja        = 0x1000da6
	sinh_tta        = 0x1000da7
	sinh_ttha       = 0x1000da8
	sinh_dda        = 0x1000da9
	sinh_ddha       = 0x1000daa
	sinh_nna        = 0x1000dab
	sinh_ndda       = 0x1000dac
	sinh_tha        = 0x1000dad
	sinh_thha       = 0x1000dae
	sinh_dha        = 0x1000daf
	sinh_dhha       = 0x1000db0
	sinh_na         = 0x1000db1
	sinh_ndha       = 0x1000db3
	sinh_pa         = 0x1000db4
	sinh_pha        = 0x1000db5
	sinh_ba         = 0x1000db6
	sinh_bha        = 0x1000db7
	sinh_ma         = 0x1000db8
	sinh_mba        = 0x1000db9
	sinh_ya         = 0x1000dba
	sinh_ra         = 0x1000dbb
	sinh_la         = 0x1000dbd
	sinh_va         = 0x1000dc0
	sinh_sha        = 0x1000dc1
	sinh_ssha       = 0x1000dc2
	sinh_sa         = 0x1000dc3
	sinh_ha         = 0x1000dc4
	sinh_lla        = 0x1000dc5
	sinh_fa         = 0x1000dc6
	sinh_al         = 0x1000dca
	sinh_aa2        = 0x1000dcf
	sinh_ae2        = 0x1000dd0
	sinh_aee2       = 0x1000dd1
	sinh_i2         = 0x1000dd2
	sinh_ii2        = 0x1000dd3
	sinh_u2         = 0x1000dd4
	sinh_uu2        = 0x1000dd6
	sinh_ru2        = 0x1000dd8
	sinh_e2         = 0x1000dd9
	sinh_ee2        = 0x1000dda
	sinh_ai2        = 0x1000ddb
	sinh_o2         = 0x1000ddc
	sinh_oo2        = 0x1000ddd
	sinh_au2        = 0x1000dde
	sinh_lu2        = 0x1000ddf
	sinh_ruu2       = 0x1000df2
	sinh_luu2       = 0x1000df3
	sinh_kunddaliya = 0x1000df4

	xf86modelock = 0x1008ff01

	xf86monbrightnessup    = 0x1008ff02
	xf86monbrightnessdown  = 0x1008ff03
	xf86kbdlightonoff      = 0x1008ff04
	xf86kbdbrightnessup    = 0x1008ff05
	xf86kbdbrightnessdown  = 0x1008ff06
	xf86monbrightnesscycle = 0x1008ff07

	xf86standby          = 0x1008ff10
	xf86audiolowervolume = 0x1008ff11
	xf86audiomute        = 0x1008ff12
	xf86audioraisevolume = 0x1008ff13
	xf86audioplay        = 0x1008ff14
	xf86audiostop        = 0x1008ff15
	xf86audioprev        = 0x1008ff16
	xf86audionext        = 0x1008ff17
	xf86homepage         = 0x1008ff18
	xf86mail             = 0x1008ff19
	xf86start            = 0x1008ff1a
	xf86search           = 0x1008ff1b
	xf86audiorecord      = 0x1008ff1c

	xf86calculator     = 0x1008ff1d
	xf86memo           = 0x1008ff1e
	xf86todolist       = 0x1008ff1f
	xf86calendar       = 0x1008ff20
	xf86powerdown      = 0x1008ff21
	xf86contrastadjust = 0x1008ff22
	xf86rockerup       = 0x1008ff23
	xf86rockerdown     = 0x1008ff24
	xf86rockerenter    = 0x1008ff25

	xf86back             = 0x1008ff26
	xf86forward          = 0x1008ff27
	xf86stop             = 0x1008ff28
	xf86refresh          = 0x1008ff29
	xf86poweroff         = 0x1008ff2a
	xf86wakeup           = 0x1008ff2b
	xf86eject            = 0x1008ff2c
	xf86screensaver      = 0x1008ff2d
	xf86www              = 0x1008ff2e
	xf86sleep            = 0x1008ff2f
	xf86favorites        = 0x1008ff30
	xf86audiopause       = 0x1008ff31
	xf86audiomedia       = 0x1008ff32
	xf86mycomputer       = 0x1008ff33
	xf86vendorhome       = 0x1008ff34
	xf86lightbulb        = 0x1008ff35
	xf86shop             = 0x1008ff36
	xf86history          = 0x1008ff37
	xf86openurl          = 0x1008ff38
	xf86addfavorite      = 0x1008ff39
	xf86hotlinks         = 0x1008ff3a
	xf86brightnessadjust = 0x1008ff3b
	xf86finance          = 0x1008ff3c
	xf86community        = 0x1008ff3d
	xf86audiorewind      = 0x1008ff3e
	xf86backforward      = 0x1008ff3f
	xf86launch0          = 0x1008ff40
	xf86launch1          = 0x1008ff41
	xf86launch2          = 0x1008ff42
	xf86launch3          = 0x1008ff43
	xf86launch4          = 0x1008ff44
	xf86launch5          = 0x1008ff45
	xf86launch6          = 0x1008ff46
	xf86launch7          = 0x1008ff47
	xf86launch8          = 0x1008ff48
	xf86launch9          = 0x1008ff49
	xf86launcha          = 0x1008ff4a
	xf86launchb          = 0x1008ff4b
	xf86launchc          = 0x1008ff4c
	xf86launchd          = 0x1008ff4d
	xf86launche          = 0x1008ff4e
	xf86launchf          = 0x1008ff4f

	xf86applicationleft  = 0x1008ff50
	xf86applicationright = 0x1008ff51
	xf86book             = 0x1008ff52
	xf86cd               = 0x1008ff53
	xf86calculater       = 0x1008ff54
	xf86clear            = 0x1008ff55
	xf86close            = 0x1008ff56
	xf86copy             = 0x1008ff57
	xf86cut              = 0x1008ff58
	xf86display          = 0x1008ff59
	xf86dos              = 0x1008ff5a
	xf86documents        = 0x1008ff5b
	xf86excel            = 0x1008ff5c
	xf86explorer         = 0x1008ff5d
	xf86game             = 0x1008ff5e
	xf86go               = 0x1008ff5f
	xf86itouch           = 0x1008ff60
	xf86logoff           = 0x1008ff61
	xf86market           = 0x1008ff62
	xf86meeting          = 0x1008ff63
	xf86menukb           = 0x1008ff65
	xf86menupb           = 0x1008ff66
	xf86mysites          = 0x1008ff67
	xf86new              = 0x1008ff68
	xf86news             = 0x1008ff69
	xf86officehome       = 0x1008ff6a
	xf86open             = 0x1008ff6b
	xf86option           = 0x1008ff6c
	xf86paste            = 0x1008ff6d
	xf86phone            = 0x1008ff6e
	xf86q                = 0x1008ff70
	xf86reply            = 0x1008ff72
	xf86reload           = 0x1008ff73
	xf86rotatewindows    = 0x1008ff74
	xf86rotationpb       = 0x1008ff75
	xf86rotationkb       = 0x1008ff76
	xf86save             = 0x1008ff77
	xf86scrollup         = 0x1008ff78
	xf86scrolldown       = 0x1008ff79
	xf86scrollclick      = 0x1008ff7a
	xf86send             = 0x1008ff7b
	xf86spell            = 0x1008ff7c
	xf86splitscreen      = 0x1008ff7d
	xf86support          = 0x1008ff7e
	xf86taskpane         = 0x1008ff7f
	xf86terminal         = 0x1008ff80
	xf86tools            = 0x1008ff81
	xf86travel           = 0x1008ff82
	xf86userpb           = 0x1008ff84
	xf86user1kb          = 0x1008ff85
	xf86user2kb          = 0x1008ff86
	xf86video            = 0x1008ff87
	xf86wheelbutton      = 0x1008ff88
	xf86word             = 0x1008ff89
	xf86xfer             = 0x1008ff8a
	xf86zoomin           = 0x1008ff8b
	xf86zoomout          = 0x1008ff8c

	xf86away        = 0x1008ff8d
	xf86messenger   = 0x1008ff8e
	xf86webcam      = 0x1008ff8f
	xf86mailforward = 0x1008ff90
	xf86pictures    = 0x1008ff91
	xf86music       = 0x1008ff92

	xf86battery   = 0x1008ff93
	xf86bluetooth = 0x1008ff94
	xf86wlan      = 0x1008ff95
	xf86uwb       = 0x1008ff96

	xf86audioforward    = 0x1008ff97
	xf86audiorepeat     = 0x1008ff98
	xf86audiorandomplay = 0x1008ff99
	xf86subtitle        = 0x1008ff9a
	xf86audiocycletrack = 0x1008ff9b
	xf86cycleangle      = 0x1008ff9c
	xf86frameback       = 0x1008ff9d
	xf86frameforward    = 0x1008ff9e
	xf86time            = 0x1008ff9f
	xf86select          = 0x1008ffa0
	xf86view            = 0x1008ffa1
	xf86topmenu         = 0x1008ffa2

	xf86red    = 0x1008ffa3
	xf86green  = 0x1008ffa4
	xf86yellow = 0x1008ffa5
	xf86blue   = 0x1008ffa6

	xf86suspend        = 0x1008ffa7
	xf86hibernate      = 0x1008ffa8
	xf86touchpadtoggle = 0x1008ffa9
	xf86touchpadon     = 0x1008ffb0
	xf86touchpadoff    = 0x1008ffb1

	xf86audiomicmute = 0x1008ffb2

	xf86keyboard = 0x1008ffb3

	xf86wwan   = 0x1008ffb4
	xf86rfkill = 0x1008ffb5

	xf86audiopreset = 0x1008ffb6

	xf86rotationlocktoggle = 0x1008ffb7

	xf86fullscreen = 0x1008ffb8

	xf86switch_vt_1  = 0x1008fe01
	xf86switch_vt_2  = 0x1008fe02
	xf86switch_vt_3  = 0x1008fe03
	xf86switch_vt_4  = 0x1008fe04
	xf86switch_vt_5  = 0x1008fe05
	xf86switch_vt_6  = 0x1008fe06
	xf86switch_vt_7  = 0x1008fe07
	xf86switch_vt_8  = 0x1008fe08
	xf86switch_vt_9  = 0x1008fe09
	xf86switch_vt_10 = 0x1008fe0a
	xf86switch_vt_11 = 0x1008fe0b
	xf86switch_vt_12 = 0x1008fe0c

	xf86ungrab        = 0x1008fe20
	xf86cleargrab     = 0x1008fe21
	xf86next_vmode    = 0x1008fe22
	xf86prev_vmode    = 0x1008fe23
	xf86logwindowtree = 0x1008fe24
	xf86loggrabinfo   = 0x1008fe25

	xf86brightnessauto = 0x100810f4
	xf86displayoff     = 0x100810f5

	xf86ok = 0x10081160

	xf86goto = 0x10081162

	xf86info = 0x10081166

	xf86vendorlogo = 0x10081168

	xf86mediaselectprogramguide = 0x1008116a

	xf86mediaselecthome = 0x1008116e

	xf86medialanguagemenu = 0x10081170
	xf86mediatitlemenu    = 0x10081171

	xf86audiochannelmode = 0x10081175

	xf86aspectratio          = 0x10081177
	xf86mediaselectpc        = 0x10081178
	xf86mediaselecttv        = 0x10081179
	xf86mediaselectcable     = 0x1008117a
	xf86mediaselectvcr       = 0x1008117b
	xf86mediaselectvcrplus   = 0x1008117c
	xf86mediaselectsatellite = 0x1008117d

	xf86mediaselecttape      = 0x10081180
	xf86mediaselectradio     = 0x10081181
	xf86mediaselecttuner     = 0x10081182
	xf86mediaplayer          = 0x10081183
	xf86mediaselectteletext  = 0x10081184
	xf86dvd                  = 0x10081185
	xf86mediaselectauxiliary = 0x10081186

	xf86audio = 0x10081188

	xf86channelup   = 0x10081192
	xf86channeldown = 0x10081193

	xf86mediaplayslow = 0x10081199

	xf86break = 0x1008119b

	xf86numberentrymode = 0x1008119d

	xf86videophone = 0x100811a0

	xf86zoomreset = 0x100811a4

	xf86editor = 0x100811a6

	xf86graphicseditor = 0x100811a8
	xf86presentation   = 0x100811a9
	xf86database       = 0x100811aa

	xf86voicemail   = 0x100811ac
	xf86addressbook = 0x100811ad

	xf86displaytoggle = 0x100811af
	xf86spellcheck    = 0x100811b0

	xf86contextmenu        = 0x100811b6
	xf86mediarepeat        = 0x100811b7
	xf8610channelsup       = 0x100811b8
	xf8610channelsdown     = 0x100811b9
	xf86images             = 0x100811ba
	xf86notificationcenter = 0x100811bc
	xf86pickupphone        = 0x100811bd
	xf86hangupphone        = 0x100811be
	xf86fn                 = 0x100811d0
	xf86fn_esc             = 0x100811d1
	xf86fnrightshift       = 0x100811e5

	xf86numeric0     = 0x10081200
	xf86numeric1     = 0x10081201
	xf86numeric2     = 0x10081202
	xf86numeric3     = 0x10081203
	xf86numeric4     = 0x10081204
	xf86numeric5     = 0x10081205
	xf86numeric6     = 0x10081206
	xf86numeric7     = 0x10081207
	xf86numeric8     = 0x10081208
	xf86numeric9     = 0x10081209
	xf86numericstar  = 0x1008120a
	xf86numericpound = 0x1008120b
	xf86numerica     = 0x1008120c
	xf86numericb     = 0x1008120d
	xf86numericc     = 0x1008120e
	xf86numericd     = 0x1008120f
	xf86camerafocus  = 0x10081210
	xf86wpsbutton    = 0x10081211

	xf86camerazoomin    = 0x10081215
	xf86camerazoomout   = 0x10081216
	xf86cameraup        = 0x10081217
	xf86cameradown      = 0x10081218
	xf86cameraleft      = 0x10081219
	xf86cameraright     = 0x1008121a
	xf86attendanton     = 0x1008121b
	xf86attendantoff    = 0x1008121c
	xf86attendanttoggle = 0x1008121d
	xf86lightstoggle    = 0x1008121e
	xf86alstoggle       = 0x10081230

	xf86refreshratetoggle = 0x10081232
	xf86buttonconfig      = 0x10081240
	xf86taskmanager       = 0x10081241
	xf86journal           = 0x10081242
	xf86controlpanel      = 0x10081243
	xf86appselect         = 0x10081244
	xf86screensaver_2     = 0x10081245
	xf86voicecommand      = 0x10081246
	xf86assistant         = 0x10081247

	xf86emojipicker             = 0x10081249
	xf86dictate                 = 0x1008124a
	xf86cameraaccessenable      = 0x1008124b
	xf86cameraaccessdisable     = 0x1008124c
	xf86cameraaccesstoggle      = 0x1008124d
	xf86accessibility           = 0x1008124e
	xf86donotdisturb            = 0x1008124f
	xf86brightnessmin           = 0x10081250
	xf86brightnessmax           = 0x10081251
	xf86kbdinputassistprev      = 0x10081260
	xf86kbdinputassistnext      = 0x10081261
	xf86kbdinputassistprevgroup = 0x10081262
	xf86kbdinputassistnextgroup = 0x10081263
	xf86kbdinputassistaccept    = 0x10081264
	xf86kbdinputassistcancel    = 0x10081265
	xf86rightup                 = 0x10081266
	xf86rightdown               = 0x10081267
	xf86leftup                  = 0x10081268
	xf86leftdown                = 0x10081269
	xf86rootmenu                = 0x1008126a
	xf86mediatopmenu            = 0x1008126b
	xf86numeric11               = 0x1008126c
	xf86numeric12               = 0x1008126d
	xf86audiodesc               = 0x1008126e
	xf863dmode                  = 0x1008126f
	xf86nextfavorite            = 0x10081270
	xf86stoprecord              = 0x10081271
	xf86pauserecord             = 0x10081272
	xf86vod                     = 0x10081273
	xf86unmute                  = 0x10081274
	xf86fastreverse             = 0x10081275
	xf86slowreverse             = 0x10081276
	xf86data                    = 0x10081277
	xf86onscreenkeyboard        = 0x10081278
	xf86privacyscreentoggle     = 0x10081279
	xf86selectivescreenshot     = 0x1008127a
	xf86nextelement             = 0x1008127b
	xf86previouselement         = 0x1008127c
	xf86autopilotengagetoggle   = 0x1008127d
	xf86markwaypoint            = 0x1008127e
	xf86sos                     = 0x1008127f
	xf86navchart                = 0x10081280
	xf86fishingchart            = 0x10081281
	xf86singlerangeradar        = 0x10081282
	xf86dualrangeradar          = 0x10081283
	xf86radaroverlay            = 0x10081284
	xf86traditionalsonar        = 0x10081285
	xf86clearvusonar            = 0x10081286
	xf86sidevusonar             = 0x10081287
	xf86navinfo                 = 0x10081288

	xf86macro1           = 0x10081290
	xf86macro2           = 0x10081291
	xf86macro3           = 0x10081292
	xf86macro4           = 0x10081293
	xf86macro5           = 0x10081294
	xf86macro6           = 0x10081295
	xf86macro7           = 0x10081296
	xf86macro8           = 0x10081297
	xf86macro9           = 0x10081298
	xf86macro10          = 0x10081299
	xf86macro11          = 0x1008129a
	xf86macro12          = 0x1008129b
	xf86macro13          = 0x1008129c
	xf86macro14          = 0x1008129d
	xf86macro15          = 0x1008129e
	xf86macro16          = 0x1008129f
	xf86macro17          = 0x100812a0
	xf86macro18          = 0x100812a1
	xf86macro19          = 0x100812a2
	xf86macro20          = 0x100812a3
	xf86macro21          = 0x100812a4
	xf86macro22          = 0x100812a5
	xf86macro23          = 0x100812a6
	xf86macro24          = 0x100812a7
	xf86macro25          = 0x100812a8
	xf86macro26          = 0x100812a9
	xf86macro27          = 0x100812aa
	xf86macro28          = 0x100812ab
	xf86macro29          = 0x100812ac
	xf86macro30          = 0x100812ad
	xf86macrorecordstart = 0x100812b0
	xf86macrorecordstop  = 0x100812b1
	xf86macropresetcycle = 0x100812b2
	xf86macropreset1     = 0x100812b3
	xf86macropreset2     = 0x100812b4
	xf86macropreset3     = 0x100812b5
	xf86kbdlcdmenu1      = 0x100812b8
	xf86kbdlcdmenu2      = 0x100812b9
	xf86kbdlcdmenu3      = 0x100812ba
	xf86kbdlcdmenu4      = 0x100812bb
	xf86kbdlcdmenu5      = 0x100812bc

	hpclearline        = 0x1000ff6f
	hpinsertline       = 0x1000ff70
	hpdeleteline       = 0x1000ff71
	hpinsertchar       = 0x1000ff72
	hpdeletechar       = 0x1000ff73
	hpbacktab          = 0x1000ff74
	hpkp_backtab       = 0x1000ff75
	hpmodelock1        = 0x1000ff48
	hpmodelock2        = 0x1000ff49
	hpreset            = 0x1000ff6c
	hpsystem           = 0x1000ff6d
	hpuser             = 0x1000ff6e
	hpmute_acute       = 0x100000a8
	hpmute_grave       = 0x100000a9
	hpmute_asciicircum = 0x100000aa
	hpmute_diaeresis   = 0x100000ab
	hpmute_asciitilde  = 0x100000ac
	hplira             = 0x100000af
	hpguilder          = 0x100000be
	hpydiaeresis       = 0x100000ee
	hplongminus        = 0x100000f6
	hpblock            = 0x100000fc

	osfcopy         = 0x1004ff02
	osfcut          = 0x1004ff03
	osfpaste        = 0x1004ff04
	osfbacktab      = 0x1004ff07
	osfbackspace    = 0x1004ff08
	osfclear        = 0x1004ff0b
	osfescape       = 0x1004ff1b
	osfaddmode      = 0x1004ff31
	osfprimarypaste = 0x1004ff32
	osfquickpaste   = 0x1004ff33
	osfpageleft     = 0x1004ff40
	osfpageup       = 0x1004ff41
	osfpagedown     = 0x1004ff42
	osfpageright    = 0x1004ff43
	osfactivate     = 0x1004ff44
	osfmenubar      = 0x1004ff45
	osfleft         = 0x1004ff51
	osfup           = 0x1004ff52
	osfright        = 0x1004ff53
	osfdown         = 0x1004ff54
	osfendline      = 0x1004ff57
	osfbeginline    = 0x1004ff58
	osfenddata      = 0x1004ff59
	osfbegindata    = 0x1004ff5a
	osfprevmenu     = 0x1004ff5b
	osfnextmenu     = 0x1004ff5c
	osfprevfield    = 0x1004ff5d
	osfnextfield    = 0x1004ff5e
	osfselect       = 0x1004ff60
	osfinsert       = 0x1004ff63
	osfundo         = 0x1004ff65
	osfmenu         = 0x1004ff67
	osfcancel       = 0x1004ff69
	osfhelp         = 0x1004ff6a
	osfselectall    = 0x1004ff71
	osfdeselectall  = 0x1004ff72
	osfreselect     = 0x1004ff73
	osfextend       = 0x1004ff74
	osfrestore      = 0x1004ff78
	osfdelete       = 0x1004ffff
}
